// 0316025 賴文揚 0316041 繆穩慶
//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      0316025 賴文揚
//----------------------------------------------
//Date:        2016/4/23
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
    );
               
//I/O ports
input   signed[16-1:0] data_i;
output  signed[32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;
always@(*)begin
	data_o <= data_i;
end

//Sign extended
          
endmodule      
     